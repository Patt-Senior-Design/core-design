../behavioral/buscmd.vh