// request defines
`define CMD_BUSRD    0
`define CMD_BUSRDX   1
`define CMD_BUSUPGR  2
`define CMD_FLUSH    3

// response defines
`define CMD_FILL     4
`define CMD_FLUSHOPT 5

// busid defines
`define BUSID_L2   0
`define BUSID_BFS  1
`define BUSID_DRAM 2
